module sine (
    input           clock, 
    input   [12:0]  p1,
    input           reset,
    output reg [9:0]  my_sine_out,
    output reg [9:0]  my_cosine_out
);

    reg [8:0] index, index_next, index_cosine;
    reg signed [9:0]LUT[511:0];
    

	always @(*)begin
        index_next = index + p1;
	end

    assign index_cosine = index+128;
	always @(posedge clock) begin
		if(reset)begin
            index   <= 0;
		end
		else begin
            index   <= index_next;
		end
    end
    assign my_sine_out = LUT[index];
    
    assign my_cosine_out = LUT[index_cosine];

    always @(posedge clock) begin
        LUT[0] <= 000;
        LUT[1] <= 006;
        LUT[2] <= 013;
        LUT[3] <= 019;
        LUT[4] <= 025;
        LUT[5] <= 031;
        LUT[6] <= 038;
        LUT[7] <= 044;
        LUT[8] <= 050;
        LUT[9] <= 056;
        LUT[10] <= 063;
        LUT[11] <= 069;
        LUT[12] <= 075;
        LUT[13] <= 081;
        LUT[14] <= 088;
        LUT[15] <= 094;
        LUT[16] <= 100;
        LUT[17] <= 106;
        LUT[18] <= 112;
        LUT[19] <= 118;
        LUT[20] <= 124;
        LUT[21] <= 130;
        LUT[22] <= 137;
        LUT[23] <= 143;
        LUT[24] <= 149;
        LUT[25] <= 155;
        LUT[26] <= 161;
        LUT[27] <= 167;
        LUT[28] <= 172;
        LUT[29] <= 178;
        LUT[30] <= 184;
        LUT[31] <= 190;
        LUT[32] <= 196;
        LUT[33] <= 202;
        LUT[34] <= 207;
        LUT[35] <= 213;
        LUT[36] <= 219;
        LUT[37] <= 225;
        LUT[38] <= 230;
        LUT[39] <= 236;
        LUT[40] <= 241;
        LUT[41] <= 247;
        LUT[42] <= 252;
        LUT[43] <= 258;
        LUT[44] <= 263;
        LUT[45] <= 269;
        LUT[46] <= 274;
        LUT[47] <= 279;
        LUT[48] <= 284;
        LUT[49] <= 290;
        LUT[50] <= 295;
        LUT[51] <= 300;
        LUT[52] <= 305;
        LUT[53] <= 310;
        LUT[54] <= 315;
        LUT[55] <= 320;
        LUT[56] <= 325;
        LUT[57] <= 330;
        LUT[58] <= 334;
        LUT[59] <= 339;
        LUT[60] <= 344;
        LUT[61] <= 348;
        LUT[62] <= 353;
        LUT[63] <= 358;
        LUT[64] <= 362;
        LUT[65] <= 366;
        LUT[66] <= 371;
        LUT[67] <= 375;
        LUT[68] <= 379;
        LUT[69] <= 384;
        LUT[70] <= 388;
        LUT[71] <= 392;
        LUT[72] <= 396;
        LUT[73] <= 400;
        LUT[74] <= 404;
        LUT[75] <= 407;
        LUT[76] <= 411;
        LUT[77] <= 415;
        LUT[78] <= 419;
        LUT[79] <= 422;
        LUT[80] <= 426;
        LUT[81] <= 429;
        LUT[82] <= 433;
        LUT[83] <= 436;
        LUT[84] <= 439;
        LUT[85] <= 442;
        LUT[86] <= 445;
        LUT[87] <= 449;
        LUT[88] <= 452;
        LUT[89] <= 454;
        LUT[90] <= 457;
        LUT[91] <= 460;
        LUT[92] <= 463;
        LUT[93] <= 465;
        LUT[94] <= 468;
        LUT[95] <= 471;
        LUT[96] <= 473;
        LUT[97] <= 475;
        LUT[98] <= 478;
        LUT[99] <= 480;
        LUT[100] <= 482;
        LUT[101] <= 484;
        LUT[102] <= 486;
        LUT[103] <= 488;
        LUT[104] <= 490;
        LUT[105] <= 492;
        LUT[106] <= 493;
        LUT[107] <= 495;
        LUT[108] <= 497;
        LUT[109] <= 498;
        LUT[110] <= 500;
        LUT[111] <= 501;
        LUT[112] <= 502;
        LUT[113] <= 503;
        LUT[114] <= 504;
        LUT[115] <= 505;
        LUT[116] <= 506;
        LUT[117] <= 507;
        LUT[118] <= 508;
        LUT[119] <= 509;
        LUT[120] <= 510;
        LUT[121] <= 510;
        LUT[122] <= 511;
        LUT[123] <= 511;
        LUT[124] <= 511;
        LUT[125] <= 511;
        LUT[126] <= 511;
        LUT[127] <= 511;
        LUT[128] <= 511;
        LUT[129] <= 511;
        LUT[130] <= 511;
        LUT[131] <= 511;
        LUT[132] <= 511;
        LUT[133] <= 511;
        LUT[134] <= 511;
        LUT[135] <= 510;
        LUT[136] <= 510;
        LUT[137] <= 509;
        LUT[138] <= 508;
        LUT[139] <= 507;
        LUT[140] <= 506;
        LUT[141] <= 505;
        LUT[142] <= 504;
        LUT[143] <= 503;
        LUT[144] <= 502;
        LUT[145] <= 501;
        LUT[146] <= 500;
        LUT[147] <= 498;
        LUT[148] <= 497;
        LUT[149] <= 495;
        LUT[150] <= 493;
        LUT[151] <= 492;
        LUT[152] <= 490;
        LUT[153] <= 488;
        LUT[154] <= 486;
        LUT[155] <= 484;
        LUT[156] <= 482;
        LUT[157] <= 480;
        LUT[158] <= 478;
        LUT[159] <= 475;
        LUT[160] <= 473;
        LUT[161] <= 471;
        LUT[162] <= 468;
        LUT[163] <= 465;
        LUT[164] <= 463;
        LUT[165] <= 460;
        LUT[166] <= 457;
        LUT[167] <= 454;
        LUT[168] <= 452;
        LUT[169] <= 449;
        LUT[170] <= 445;
        LUT[171] <= 442;
        LUT[172] <= 439;
        LUT[173] <= 436;
        LUT[174] <= 433;
        LUT[175] <= 429;
        LUT[176] <= 426;
        LUT[177] <= 422;
        LUT[178] <= 419;
        LUT[179] <= 415;
        LUT[180] <= 411;
        LUT[181] <= 407;
        LUT[182] <= 404;
        LUT[183] <= 400;
        LUT[184] <= 396;
        LUT[185] <= 392;
        LUT[186] <= 388;
        LUT[187] <= 384;
        LUT[188] <= 379;
        LUT[189] <= 375;
        LUT[190] <= 371;
        LUT[191] <= 366;
        LUT[192] <= 362;
        LUT[193] <= 358;
        LUT[194] <= 353;
        LUT[195] <= 348;
        LUT[196] <= 344;
        LUT[197] <= 339;
        LUT[198] <= 334;
        LUT[199] <= 330;
        LUT[200] <= 325;
        LUT[201] <= 320;
        LUT[202] <= 315;
        LUT[203] <= 310;
        LUT[204] <= 305;
        LUT[205] <= 300;
        LUT[206] <= 295;
        LUT[207] <= 290;
        LUT[208] <= 284;
        LUT[209] <= 279;
        LUT[210] <= 274;
        LUT[211] <= 269;
        LUT[212] <= 263;
        LUT[213] <= 258;
        LUT[214] <= 252;
        LUT[215] <= 247;
        LUT[216] <= 241;
        LUT[217] <= 236;
        LUT[218] <= 230;
        LUT[219] <= 225;
        LUT[220] <= 219;
        LUT[221] <= 213;
        LUT[222] <= 207;
        LUT[223] <= 202;
        LUT[224] <= 196;
        LUT[225] <= 190;
        LUT[226] <= 184;
        LUT[227] <= 178;
        LUT[228] <= 172;
        LUT[229] <= 167;
        LUT[230] <= 161;
        LUT[231] <= 155;
        LUT[232] <= 149;
        LUT[233] <= 143;
        LUT[234] <= 137;
        LUT[235] <= 130;
        LUT[236] <= 124;
        LUT[237] <= 118;
        LUT[238] <= 112;
        LUT[239] <= 106;
        LUT[240] <= 100;
        LUT[241] <= 094;
        LUT[242] <= 088;
        LUT[243] <= 081;
        LUT[244] <= 075;
        LUT[245] <= 069;
        LUT[246] <= 063;
        LUT[247] <= 056;
        LUT[248] <= 050;
        LUT[249] <= 044;
        LUT[250] <= 038;
        LUT[251] <= 031;
        LUT[252] <= 025;
        LUT[253] <= 019;
        LUT[254] <= 013;
        LUT[255] <= 006;
        LUT[256] <= 000;
        LUT[257] <= -06;
        LUT[258] <= -13;
        LUT[259] <= -19;
        LUT[260] <= -25;
        LUT[261] <= -31;
        LUT[262] <= -38;
        LUT[263] <= -44;
        LUT[264] <= -50;
        LUT[265] <= -56;
        LUT[266] <= -63;
        LUT[267] <= -69;
        LUT[268] <= -75;
        LUT[269] <= -81;
        LUT[270] <= -88;
        LUT[271] <= -94;
        LUT[272] <= -100;
        LUT[273] <= -106;
        LUT[274] <= -112;
        LUT[275] <= -118;
        LUT[276] <= -124;
        LUT[277] <= -130;
        LUT[278] <= -137;
        LUT[279] <= -143;
        LUT[280] <= -149;
        LUT[281] <= -155;
        LUT[282] <= -161;
        LUT[283] <= -167;
        LUT[284] <= -172;
        LUT[285] <= -178;
        LUT[286] <= -184;
        LUT[287] <= -190;
        LUT[288] <= -196;
        LUT[289] <= -202;
        LUT[290] <= -207;
        LUT[291] <= -213;
        LUT[292] <= -219;
        LUT[293] <= -225;
        LUT[294] <= -230;
        LUT[295] <= -236;
        LUT[296] <= -241;
        LUT[297] <= -247;
        LUT[298] <= -252;
        LUT[299] <= -258;
        LUT[300] <= -263;
        LUT[301] <= -269;
        LUT[302] <= -274;
        LUT[303] <= -279;
        LUT[304] <= -284;
        LUT[305] <= -290;
        LUT[306] <= -295;
        LUT[307] <= -300;
        LUT[308] <= -305;
        LUT[309] <= -310;
        LUT[310] <= -315;
        LUT[311] <= -320;
        LUT[312] <= -325;
        LUT[313] <= -330;
        LUT[314] <= -334;
        LUT[315] <= -339;
        LUT[316] <= -344;
        LUT[317] <= -348;
        LUT[318] <= -353;
        LUT[319] <= -358;
        LUT[320] <= -362;
        LUT[321] <= -366;
        LUT[322] <= -371;
        LUT[323] <= -375;
        LUT[324] <= -379;
        LUT[325] <= -384;
        LUT[326] <= -388;
        LUT[327] <= -392;
        LUT[328] <= -396;
        LUT[329] <= -400;
        LUT[330] <= -404;
        LUT[331] <= -407;
        LUT[332] <= -411;
        LUT[333] <= -415;
        LUT[334] <= -419;
        LUT[335] <= -422;
        LUT[336] <= -426;
        LUT[337] <= -429;
        LUT[338] <= -433;
        LUT[339] <= -436;
        LUT[340] <= -439;
        LUT[341] <= -442;
        LUT[342] <= -445;
        LUT[343] <= -449;
        LUT[344] <= -452;
        LUT[345] <= -454;
        LUT[346] <= -457;
        LUT[347] <= -460;
        LUT[348] <= -463;
        LUT[349] <= -465;
        LUT[350] <= -468;
        LUT[351] <= -471;
        LUT[352] <= -473;
        LUT[353] <= -475;
        LUT[354] <= -478;
        LUT[355] <= -480;
        LUT[356] <= -482;
        LUT[357] <= -484;
        LUT[358] <= -486;
        LUT[359] <= -488;
        LUT[360] <= -490;
        LUT[361] <= -492;
        LUT[362] <= -493;
        LUT[363] <= -495;
        LUT[364] <= -497;
        LUT[365] <= -498;
        LUT[366] <= -500;
        LUT[367] <= -501;
        LUT[368] <= -502;
        LUT[369] <= -503;
        LUT[370] <= -504;
        LUT[371] <= -505;
        LUT[372] <= -506;
        LUT[373] <= -507;
        LUT[374] <= -508;
        LUT[375] <= -509;
        LUT[376] <= -510;
        LUT[377] <= -510;
        LUT[378] <= -511;
        LUT[379] <= -511;
        LUT[380] <= -511;
        LUT[381] <= -512;
        LUT[382] <= -512;
        LUT[383] <= -512;
        LUT[384] <= -512;
        LUT[385] <= -512;
        LUT[386] <= -512;
        LUT[387] <= -512;
        LUT[388] <= -511;
        LUT[389] <= -511;
        LUT[390] <= -511;
        LUT[391] <= -510;
        LUT[392] <= -510;
        LUT[393] <= -509;
        LUT[394] <= -508;
        LUT[395] <= -507;
        LUT[396] <= -506;
        LUT[397] <= -505;
        LUT[398] <= -504;
        LUT[399] <= -503;
        LUT[400] <= -502;
        LUT[401] <= -501;
        LUT[402] <= -500;
        LUT[403] <= -498;
        LUT[404] <= -497;
        LUT[405] <= -495;
        LUT[406] <= -493;
        LUT[407] <= -492;
        LUT[408] <= -490;
        LUT[409] <= -488;
        LUT[410] <= -486;
        LUT[411] <= -484;
        LUT[412] <= -482;
        LUT[413] <= -480;
        LUT[414] <= -478;
        LUT[415] <= -475;
        LUT[416] <= -473;
        LUT[417] <= -471;
        LUT[418] <= -468;
        LUT[419] <= -465;
        LUT[420] <= -463;
        LUT[421] <= -460;
        LUT[422] <= -457;
        LUT[423] <= -454;
        LUT[424] <= -452;
        LUT[425] <= -449;
        LUT[426] <= -445;
        LUT[427] <= -442;
        LUT[428] <= -439;
        LUT[429] <= -436;
        LUT[430] <= -433;
        LUT[431] <= -429;
        LUT[432] <= -426;
        LUT[433] <= -422;
        LUT[434] <= -419;
        LUT[435] <= -415;
        LUT[436] <= -411;
        LUT[437] <= -407;
        LUT[438] <= -404;
        LUT[439] <= -400;
        LUT[440] <= -396;
        LUT[441] <= -392;
        LUT[442] <= -388;
        LUT[443] <= -384;
        LUT[444] <= -379;
        LUT[445] <= -375;
        LUT[446] <= -371;
        LUT[447] <= -366;
        LUT[448] <= -362;
        LUT[449] <= -358;
        LUT[450] <= -353;
        LUT[451] <= -348;
        LUT[452] <= -344;
        LUT[453] <= -339;
        LUT[454] <= -334;
        LUT[455] <= -330;
        LUT[456] <= -325;
        LUT[457] <= -320;
        LUT[458] <= -315;
        LUT[459] <= -310;
        LUT[460] <= -305;
        LUT[461] <= -300;
        LUT[462] <= -295;
        LUT[463] <= -290;
        LUT[464] <= -284;
        LUT[465] <= -279;
        LUT[466] <= -274;
        LUT[467] <= -269;
        LUT[468] <= -263;
        LUT[469] <= -258;
        LUT[470] <= -252;
        LUT[471] <= -247;
        LUT[472] <= -241;
        LUT[473] <= -236;
        LUT[474] <= -230;
        LUT[475] <= -225;
        LUT[476] <= -219;
        LUT[477] <= -213;
        LUT[478] <= -207;
        LUT[479] <= -202;
        LUT[480] <= -196;
        LUT[481] <= -190;
        LUT[482] <= -184;
        LUT[483] <= -178;
        LUT[484] <= -172;
        LUT[485] <= -167;
        LUT[486] <= -161;
        LUT[487] <= -155;
        LUT[488] <= -149;
        LUT[489] <= -143;
        LUT[490] <= -137;
        LUT[491] <= -130;
        LUT[492] <= -124;
        LUT[493] <= -118;
        LUT[494] <= -112;
        LUT[495] <= -106;
        LUT[496] <= -100;
        LUT[497] <= -94;
        LUT[498] <= -88;
        LUT[499] <= -81;
        LUT[500] <= -75;
        LUT[501] <= -69;
        LUT[502] <= -63;
        LUT[503] <= -56;
        LUT[504] <= -50;
        LUT[505] <= -44;
        LUT[506] <= -38;
        LUT[507] <= -31;
        LUT[508] <= -25;
        LUT[509] <= -19;
        LUT[510] <= -13;
        LUT[511] <= -06;

    end
    endmodule